PK   繞W�e��,#  LY    cirkitFile.json�ݎ�F��_��b�d&���c쌍�`���A�b�-Lu�W���6���e��6���J�(�'�vz�q��<�L����]�c����]�~����~�����]�k��jnV6��~[���?�[����N��|I�u�lc�ʇ2t�	I��6q뚒�f!I�u���vEg���ի�oo^�@b��!f�*�ʊ�
�J�RS91�T�T^� U0U&f�*�*3HLU��
�*�R��!O�b�(H��\I�d)��"�t)��"�)��"�)��"�)��"�)��"��)��"���>l
�dWo��T�w�n��%�?��{$��V��{�'������}��W67�Bl�ĥ�I�uf��M�ufm\T�{ ��b�H��s���p�D���p�D���p�D���p�D���p�D���p�D����2`�]>l�0���T��c��<��/�+�y��%$�*���ET�>�_KR��D,)���D��_K��B~-KD
��D,)������<��%"	�WL�@o��cz'��Ί�J�0�;yKD
�Mpyw�.���.���.���.���.�0���p�D������B�w��B�;��B�;���Q�;�<w�%"�<w�%"�<w�%"�<w�%L��s�X"R�s�X"R�s�Hb�Pޜ��ʱ1�����t,�ac�#,��,6v;(a�L�bc�bc�#,]���9l�t���cl�����ݗڬ�҇<q�7���4)Z
I�4�)K�_��,N�����aÞa�,���t�ʱ�˱�����T6v6vP:�ҙ��Ʈ��JGX:�p
W�M	���|<U?�1A;�5!�7!�9�����'��6(X>���jp��&�G`>��t<O`>��dvp����G`>����u`�����;,��NW.@�7�K{P)�Y��=:�{�[�`�b���G`>^%�ؾ`����[��C?[A?\��/l_�|��5E�������|�
?�}�����q���/X>��
4p����G`>^;�ؾ`��7^q'����2H�����K��K���G`>^ 	�ؾ`��w�4��=����
�^`w���0\��e��e��e`����O
v?X>���]p����G`>^y���`���k����,��x�78~`���#0�S�l_�|�����9�}����ti?$~#{ yx�H8�����=a���ǁ�`���e���,��� 8~�2�2`����Ł����|\t?�}����˅���/X>�q�p����G`>.��ؾ`����e���`���#0������G`>.���`��ǥ����,����8~`���#0���?�|���U�������|\r?�����������X>�q�3p����G`>.І�_�X>�qi9p�.<>YX�8>:����5a�F��šr�9����w�7�[�a=ƥo�5V@\�|X�uqG�RXʰh��� ܓ%��K�.l>����������,=������K�ψ�+������k�������u/��п�M����;z����	'X�v�Z�ϓ��'��]jK�O�M��fUa��Nxލ^7�����d�G/[�~��ѵ�MC�$�(b�,͓��!���	E]��Aܬ��_��f�j~ᬳ!���N�"��ٺ�ͳ,qm�5i��� vN��}/����ubŞ�&)s�%�����2����볚O��1�Ǯb�66o�uR��E0)����&\��Yͧ}]���M3F�%.4eҸ.$�:�u�gm�.����ӿ>�j�l���xgfNɫ������v��V���v�z����p`V�b�?�IN	�$d8ea�@B�� �$d�c�@B�M2�$d�wc�@B��7�$d��c�@B�o`�@B��� J����K۰�M�čR2�=,w,y��Lo���K�(%���1�r8��8J�/E��(���	�`y����Q)�B&XG)��N�	��-,���LK�����QJ���	b��q��(%��g1���J_-gJay��Tc� d�����B&X?(ɯ�\����),�����
�	��SXG)q,���<�R�Z0&�x���8J��� �-6w�<~P���2��8J��Ø`y���8J�nØ`y���8J�Ø`y���8J�����򸇍�QJ�`����ay��aL����Ǜ�<�ay�ċ�`L�<�ay�ċ�`L�<���8J��Ø`y<���)����k���Z�*���
+�j�u�<VRa5�p�\WVRa5հ\WVRa��K%��
�h��
��D_`\��+���{��p���Yֲ����+���jX��
��+���jX��
��+���jX�
��+���`c��ThI���6��V�u)�.�E:Ƌt��
-���\s���/Zҡ�9�:��q`*��C�s�ub��lH��thy�Nlu��
-���Z���1Zҡ�5%:��qd*��C�kctb;v:��^*�t���ˬ�/S�%Z^��[_�BK:���J'�JOĔ���2��ˬ�/S�%Z^�[_�BK:���O'�:�L��thyM�Nlu|�
-����J����2Zҡ�5�:���e*��C�k]G���2Ydlu|�
-��ՙ����ThI�����VǗ�В-��։��� �ը��9ZH�&+*�VT�����R_���2Zҡ��:���e*��C�5tb���ThI��k%��VǗ�В-�|Љ��/S�%Z�]�[_�BK:�\�C%�NǗ�В-�щ��� ��
-���AǗ9��e*��C˵]tb���ThI��k���Vi%��R2_�t|���e*��C�5�tb���ThI��k��VǗ�В-�p҉��/S�%Z�E�[_�BK:�\SK%�^Ǘ�В-�Ӊ���2Zҡ�g:���e*��C˵�tb���ThI��k���VǗ�В-��Ӊ��/S�%Z��[_�BK:�\�P'�:�L��th�&�Nlu|�
-��rmI����2Zҡ��*��t|�
-��r�O���</S��s�� ��bns����Тe'i�"z���B��ڴK_WQ���Pŝ�bU&je/T�Ο�U&�Q/T�� �Pe����^꼘�;��ץ2��;�jե2�<�ӥ2�>||M����Ke0�x굞Ke�^<~�R�C/��m��O�Xr�����Fߥ�DӋ�^��T����w*-��bz��{�d�6�ih�$E���<ih�ڛΘP�uQ_��R��\�,�R�~>��YW'e�Q�l�E�,K\۬CAM��1ڛ�r5.�q�X�Nl�8��]�������MLRuy�e��Uc��=+ĶmTi�uR��[E0)����&\g��r�e]���M��.��2i\c��ȳ�u�Yf�\e��:+}ȣ�7���4)ڸ�EӬӦ,}f�����s�
=K��z�j����>�^}|�]�*���]}��o��,@B��WH���B2}.���L�� D !�;GH��.B2�����L�!D !�;mH�\;&E�6.m��6�7J�nN`�`��`��d�M0L��M��R2�:&X'XG)�í&,�[XG)��M0n������q��9���0���q��9܅�0���q��9��0���q��9ܹ��qXOay��5�`L�;)�[)�<���8J�k���`y<��q��B�1��x
��(%��c��q��(%�� c��q��(%�- c������q��(%^c��q��(%^sc��q��(%^�
{�����QJ�������QJ��Ƅ{��{�	����QJ��
�����QJ�����,���x-	�	��3X�RZ�.d���zX�P%VRae]����A"��J*���7B���J*��Հ@���J*��w��uT�VRa�� ���J?@"��J*�q���Q�H4XI��T��hU`\5XI��T�zhU`\5XI��T�ZhU`\5XI����ǥBK:�<�Y'�J�K�v��.�1^��ThI�����V�}�В-ϙ׉��S�%Z���[�BK:���A'�:NL��thy-�Nluܘ
-������82Zҡ�1:��qe*��C�k|t,��2Zҡ�J:���e*��C�k�tb��DL鑘�/�:����2Zҡ�5p:���e*��C�k�tb���ThI���$��VǗ�В-��ԉ��/S�%Z^#�[_�BK:���U'�:�L��thyͮ��$_�BK:���X'�:�L��thy�Nlu|�
-���Zp��*�VT�����R_���2Zҡ��:���e*��C�5tb���ThI��k%��VǗ�В-�|Љ��/S�%Z�]�[_�BK:�\�C%�NǗ�В-�щ��/S�%Z���[_�BK:�\�E'�:�L��th�F�Nl�V�)-%��eNǗ9_�BK:�\3H'�:�L��th���Nlu|�
-��r'����2Zҡ�ZT:���e*��C�5�Tb�u|�
-��rm0����2Zҡ�g:���e*��C˵�tb���ThI��k���VǗ�В-��Ӊ�R��2:����2���ThI��k��VǗ�В-�dԉ��/S�%Z�-�[_�BK:�\#S%���/S�%Z���[_�BK:�\�T'�:�L����.|��D�ۅ*�i�LT�]�F{��D��*���LT�^�2Q�z��D�*5���:P���ީ��.���ߩW�.�����.����ׄ.���⩗q.��`L/�zK�RL/�z�RL/�z��RL/�z��ҫ.�O�=�I�kC���IBQD�,͓��!���	E]��Q�,��j����Ɇ�κ:)��g�.�dY��f
j�������q)����ub���M�t>�o�`��:�,��,�8{V�mۨ�t��q��`R*��M��2K�*˺�m��"q]�%.4eҸ.$�:�u�gm뮳�R��R�uV��Go��iR�q��Y�MY����,�T��|���9���n��6�ϫW�f��f�w�:�����ڰ[�z���7_�o�9��y{#�q$�W@@�~�!����8+����$CI��F�Ҿ!<s�k�������O虳�{@ϔ壽����p��b�o���(��,��s����-{Fr�DY|���o����qXP߷�F�#d����}���װ	B=�Q*�X
B%Ra(�#+L�A�0�A��z���	ɒ�A�<6�����o<P��
�+�u�~�4�9�>C�ێ��@�a5������V�zV�>�{�u�j��7���Gɘ��V�y������>
)��
 �K��)��B,a��B
����f)����!�K�~n��B,a��%B
����)��0�E����>�� 	T�a�s��J�$*�0�	BR@%@"�k��%) � ��5�a���bҫ��^c�gV�ȶrs�&� d[ȶrs��&� d[ȶrs�	'� d[ȶrs��'� d[��3;�N@�M�d[/�d�^c��X���k�r!�� ��\,��z� @.N�X��ut�\�r�\��8 C]H�r��	�(%�0�u�l��d�T�ȶr��� d[ȶr��� d[ȶr�$� d[ȶr�Px� ȶ0��kp�+ �N��S�WTp �~!��S�W�p ��S�WKp �iȧr��� ���O��g��*����-Dz�#0+b�7*�"�_,��L5���Ӄ��G`>S��[�� ����/�p�F�+����#0���HH�F�)7�D9	�Kc\��
S�� ��G`>S��O�� �����T��8=H��|�3ը�$N?,��x�$z<�6$`BB�TOt��Jж�о���LHhB�b��!ڜ�		M�Ӄ�1D0!�	yj3:��Q?�		M�Ӳ�1D;0!�	yJ9:�hw&$4!O�G��P���&4'�=01��K^�kK�:�m�E�0!�	y�:�h�&$4!��@��<�@m[,ڶX�m���٠c��-`BB�!tѶLHhB^߄�!ڶ�		M�k��1D�0!�	y]:�h�&$4�V���m2}LHѶL���гGжLHhB^|��!ڶ�		MxZpÑ)����@��1�4��a�a�ah��]L�v1`BB��Zt�.LHh�q�H� &�h&�U���]��Є�"C����W��c��-`BB�Jxpڶ�		MxZGÑ)�T#�@��1�4h��_���&�r	��m��Є\�C�����mqh��жLHhB.���!ڶ�		M��A�1D�0!�	��	:�h�&$4!�eA�m[���&�2�z�m����c�~�&$4!��A��S���&�2D��}
��Є\B	C�O���?�c��)`BBr�*t�>LHhB.���!ڧ�		M�%��1D�0!�	��:�h�&$4!�j�0C�0!�	O_����+�7��� K#02�8}L/E��+��"9*��������ۏ��.~����PnTCu�kN/���F%L��]�~T2ti�wOi��en�������T@�)�oR[* �������㗎-M[Ҏiϼ?�K�μ��I���v�����nk�ɔD/\����;���M��)�^<��x�Υ'��m�&	E�4OZ����3&u]ԗ���K�Bv����YbCXg]��EF��u�gY��f
j�����ל���0�k׉���k�27]����)���K�?���ߏ���>b�6�o�uR��E0)����&\��Y�/����m��"q]�%.4eҸ.$�:�u�gm�.����~��/�6]�>�3����If������~�I�z�z�L�:���	��,|���v�����<N���$K�)��oM�9����[Xna{mna����[Xna����[��"&��7�9���-���s�al0�d8i0���4���N����^�x8��a�Ǿ�_���������7Ċ���(˘���N4u<�uL�D��UU4y)�DR�;�eB"+�g�e�c�\3+#.Zi%G5��1Q*$rS�Ę�8!��o��iӕR�A.��x���`��F���J�'���l��b�?﫻�	w|M^��9��X���W4���r���+?�*;~���ʏ_����+;�*=~���*�_���W��+�54}G?\���g�cs�m���Þ���������{U�ݖ��P�����\u�=����G?�����<^����n�!���Џ�����p���z��6�|���������������e��#<�o"�*������o��5�^u��C�_>���6��.|�l��q����>�H<���Ǯ^�waw	��f�Hv���~ �(1�n��m��k"���yg��S{�c4��*Z���ΤI�c"ȝY'��MLi�$���6�	������?t���6�p������z�[߅�|]F��"�<���O��>O�}�}�=��x�y??9�_X������?�<�yq*D��Sc�^Ħ�4�'y#~�Ӊ/���T�r��T��m�d?�&�l3����,�wv��X���?rg��m��6�c|n��o�������?����������6��1YK����sB�g�� ]}�������{�|��J3J]�������֕�;~R��y�:�M�RJ�'-��[��m^�!M����k�ݐy�˝\�nlQ.^������v�٣^q����)��8�C�qG�";n�����2����������T����n[�qw��1�消g��?vGS���柏��޸���]}�y�%yWg	��'YQ��]�z�[l3zc���&�Y��؁��fg6�g�A������O�%��<�v�Y�\gt �J��3���%��3_����%<l{�����G���l���f��2�#���38f|8���o�i�R���7��MM�L�]��Ά��ۻ��D�v�����VO@�����r{�G����������i����Lw��??�o��o�/���ۇ�|�m�(�	���7٬�����)�̷i�X��������:��س��N�B�x_�$P�9������={ֳ�a��m~x����Mjܙ�x&����g��Ե�$��>�v�YO��u�s�î}4A����f����˶�v����ܷ��&<��6��$��'��O�y~��x���غ���L��\��hb�X��I�X��6��!j'=h�c�a:�H��h��s�h�^Jd�����u	��}����~�o|z��Y?��o޽Z%i����[I?m����a����ޅ�sǳ�e�֤%���Ö�����z�.�_}���.����m~��x`�T��M�w�ݛի7�����+�fu�&��z��ns�M�%z���������n�����*o���$��?����GE������z�����͛�1�������?g��W���O/��7[x��3[ſ�z����S�4�������: OMCw�s�;@��jl5�2&ˡ��"\� �g&h���2؅����t�R����VޝߊoV/ު��Y�{6E@w�,��Y��Ћ:���t�ӭ��?�X�����������b�c��|��c���v�rN�9���p��ȂgGA�`��b���~i.Ig��ECK}�/T(����v�wpsN��V��r���|Ѹ��7�Uܥ\�x��^WqWs��`���bN.l5��^d�V�q��9�Ћ�`�絎�"V�e���ˈ?9�E>�9N�*���y+���m�,� ��:��t���u��6��j׻��V�����l�Q�t�3��������s�v�Ȧ�M��8��7g7�;x5�KKd���R�҉���`����-�9�s�U6qԟ�,�lb�u6ww�v��a���K�/�?6��?�����W������ޥ��V��PK
   繞W�e��,#  LY                  cirkitFile.jsonPK      =   Y#    